module contador ( 
	en,
	clr,
	clk,
	display
	) ;

input  en;
input  clr;
input  clk;
inout [6:0] display;
