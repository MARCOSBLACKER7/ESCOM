LIBRARY IEEE;   
USE IEEE.STD_LOGIC_1164.ALL;    
    
ENTITY TECLADO IS         
    PORT (
	   	CLK, CLR: IN STD_LOGIC;
		FILA: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		COLUMNA: INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	    D: INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
    );

    ATTRIBUTE PIN_NUMBERS OF TECLADO : ENTITY IS
	"CLK:1 "		&
	"CLR:13 "		&
	"FILA(3):11 "	&
	"FILA(2):10 "	&
	"FILA(1):9 "	&
	"FILA(0):8 "	&
    "D(0):15 "   	&   
    "D(1):16 "   	&   
    "D(2):17 "   	&  
    "D(3):18 "   	&  
	"D(4):19 "   	&  
	"D(5):20 "   	&  
	"D(6):21 "      &
 	"COLUMNA(0):14 "    &
	"COLUMNA(1):22 "    &
	"COLUMNA(2):23 ";
END TECLADO;  

ARCHITECTURE PROGRAMA OF TECLADO IS 
	CONSTANT ASTERISCO : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0001000";
	CONSTANT GATO : STD_LOGIC_VECTOR(6 DOWNTO 0):=  "0000100";
	CONSTANT CERO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0000001";
	CONSTANT UNO  :  STD_LOGIC_VECTOR(6 DOWNTO 0):=    "1001111";
	CONSTANT DOS  :  STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0010010";
	CONSTANT TRES : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0000110";
	CONSTANT CUATRO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "1001100";
	CONSTANT CINCO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0100100";
	CONSTANT SEIS : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0100000";
	CONSTANT SIETE : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0001111";
	CONSTANT OCHO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0000000";
	CONSTANT NUEVE : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0000100";
	SIGNAL L: STD_LOGIC;
	SIGNAL LLAVE: STD_LOGIC_VECTOR(6 DOWNTO 0);

	  BEGIN
	  --COMPUERTA LOGICA
			L<= NOT(FILA(0) AND FILA(1) AND FILA(2) AND FILA(3));
	  --CONTADOR DE ANILLO
			PANILLO : PROCESS(CLK,CLR)
			BEGIN
				IF(CLR = '1') THEN
					COLUMNA<="110";
				ELSIF(RISING_EDGE(CLK)) THEN
 				    COLUMNA<=TO_STDLOGICVECTOR(TO_BITVECTOR(COLUMNA) ROL 1);
				END IF;
			END PROCESS PANILLO;
	  --CONVERTIDOR DE CODIGO
			TECLA: PROCESS(FILA,COLUMNA)
			BEGIN
				CASE FILA&COLUMNA IS
				WHEN "0111101"=>
					LLAVE<= CERO;
				WHEN "1110011"=>
					LLAVE<= UNO;
				WHEN "1110101"=>
					LLAVE<= DOS;
				WHEN "1110110"=>
					LLAVE<= TRES;
				WHEN "1101011"=>
					LLAVE<= CUATRO;
			   	WHEN "1101101"=>
					LLAVE<= CINCO;
				WHEN "1101110"=>
					LLAVE<= SEIS;
				WHEN "1011011"=>
					LLAVE<= SIETE;
				WHEN "1011101"=>
					LLAVE<= OCHO;
				WHEN "1011110"=>
					LLAVE<= NUEVE;
				WHEN "0111110"=>
					LLAVE<= GATO;
				WHEN "0111011"=>
					LLAVE<= ASTERISCO;
				WHEN OTHERS=>
					LLAVE<=(OTHERS => '-');
				END CASE;
			END PROCESS TECLA;
		--REGISTRO
			REGISTRO: PROCESS(CLK,CLR)
			BEGIN
				IF(CLR = '1') THEN
					D <= (OTHERS=>'1');
				ELSIF(RISING_EDGE(CLK)) THEN
 				    CASE L IS
						WHEN '0' =>
						 D <= D;
						WHEN OTHERS =>
						 D <= LLAVE;
					END CASE;
				END IF;
			END PROCESS REGISTRO;
END PROGRAMA;