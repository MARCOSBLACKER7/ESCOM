Library IEEE;   
Use IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
   

ENTITY SENSOR IS
    PORT (CLK, CLR: IN STD_LOGIC;  
    UNI: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    DEC: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    SENSORES: IN STD_LOGIC_VECTOR(1 downto 0)
    );
ATTRIBUTE PIN_NUMBERS OF SENSOR : ENTITY IS
"CLK:1          "   &
"CLR:13         "	&
"SENSORES(0):2   "	& --SENSORES
"SENSORES(1):3   "	&
"DEC(2):20      "	& --DECENAS
"DEC(1):19      "	&
"DEC(0):18      "	&
"UNI(3):17      "	& --UNIDADES
"UNI(2):16      "	&
"UNI(1):15      "	&
"UNI(0):14      ";
END SENSOR;  

ARCHITECTURE PROGRAMA OF SENSOR IS
TYPE STATES IS (Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7);  
SIGNAL ESTADO_PRESENTE, ESTADO_SIGUIENTE: STATES; --ESTADOS
SIGNAL PCONTADOR: STD_LOGIC_VECTOR(1 downto 0);
BEGIN 
MAQUINAESTADOS : PROCESS(ESTADO_PRESENTE, SENSORES) --AUTOMATA
BEGIN
CASE ESTADO_PRESENTE IS
    WHEN Q0 => 
        CASE SENSORES IS
            WHEN "00" => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="00";
            WHEN "01" => 
ESTADO_SIGUIENTE <= Q4;
PCONTADOR <="00";
            WHEN "10" => 
ESTADO_SIGUIENTE <= Q1;
PCONTADOR <="00";
            WHEN OTHERS => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="00";
        END CASE;
WHEN Q1 => 
        CASE SENSORES IS
            WHEN "00" => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="00";
            WHEN "01" => 
ESTADO_SIGUIENTE <= Q4;
PCONTADOR <="00";
            WHEN "10" => 
ESTADO_SIGUIENTE <= Q1;
PCONTADOR <="00";
            WHEN OTHERS => 
ESTADO_SIGUIENTE <= Q2;
PCONTADOR <="00";
        END CASE;
WHEN Q2 => 
        CASE SENSORES IS
            WHEN "00" => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="00";
            WHEN "01" => 
ESTADO_SIGUIENTE <= Q3;
PCONTADOR <="00";
            WHEN "10" => 
ESTADO_SIGUIENTE <= Q1;
PCONTADOR <="00";
            WHEN OTHERS => 
ESTADO_SIGUIENTE <= Q2;
PCONTADOR <="00";
        END CASE;
WHEN Q3 => 
        CASE SENSORES IS
            WHEN "00" => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="01";
            WHEN "01" => 
ESTADO_SIGUIENTE <= Q3;
PCONTADOR <="00";
            WHEN "10" => 
ESTADO_SIGUIENTE <= Q1;
PCONTADOR <="01";
            WHEN OTHERS => 
ESTADO_SIGUIENTE <= Q2;
PCONTADOR <="00";
        END CASE;
WHEN Q4 => 
        CASE SENSORES IS
            WHEN "00" => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="00";
            WHEN "01" => 
ESTADO_SIGUIENTE <= Q4;
PCONTADOR <="00";
            WHEN "10" => 
ESTADO_SIGUIENTE <= Q1;
PCONTADOR <="00";
            WHEN OTHERS => 
ESTADO_SIGUIENTE <= Q5;
PCONTADOR <="00";
        END CASE;
WHEN Q5 => 
        CASE SENSORES IS
            WHEN "00" => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="00";
            WHEN "01" => 
ESTADO_SIGUIENTE <= Q4;
PCONTADOR <="00";
            WHEN "10" => 
ESTADO_SIGUIENTE <= Q6;
PCONTADOR <="00";
            WHEN OTHERS => 
ESTADO_SIGUIENTE <= Q5;
PCONTADOR <="00";
        END CASE;
WHEN Q6 => 
        CASE SENSORES is
            WHEN "00" => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="10";
            WHEN "01" => 
ESTADO_SIGUIENTE <= Q4;
PCONTADOR <="10";
            WHEN "10" => 
ESTADO_SIGUIENTE <= Q6;
PCONTADOR <="00";
            WHEN OTHERS => 
ESTADO_SIGUIENTE <= Q5;
PCONTADOR <="00";
        END CASE;
WHEN Q7 => 
        CASE SENSORES IS
            WHEN "00" => 
ESTADO_SIGUIENTE <= Q0;
PCONTADOR <="00";
            WHEN "01" => 
ESTADO_SIGUIENTE <= Q4;
PCONTADOR <="00";
            WHEN "10" => 
ESTADO_SIGUIENTE <= Q1;
PCONTADOR <="00";
            WHEN OTHERS => 
ESTADO_SIGUIENTE <= Q7;
PCONTADOR <="00";
        END CASE;
END CASE;
END PROCESS MAQUINAESTADOS;

PROCESS(CLK, CLR)
BEGIN
IF CLR = '1' THEN 
	ESTADO_PRESENTE <=Q0;
ELSIF RISING_EDGE(CLK) THEN
	ESTADO_PRESENTE <= ESTADO_SIGUIENTE;
END IF;
END PROCESS;

CONTADOR_DECADA: PROCESS(CLK, CLR)
BEGIN
IF CLR = '1' THEN
	UNI <= (OTHERS => '0');
	DEC <= (OTHERS => '0');
ELSIF RISING_EDGE(CLK) THEN
	IF PCONTADOR = "00" THEN
		UNI <= UNI;
		DEC <= DEC;
	END IF;

	IF PCONTADOR = "01" THEN
		UNI <= UNI + 1;

		IF UNI = "1001" THEN
			UNI <= "0000";
			DEC <= DEC + 1;
		END IF;
	END IF;

	IF PCONTADOR = "10" THEN
		UNI <= UNI - 1;

		IF UNI = "0000" THEN
			UNI <= "1001";
			DEC <= DEC - 1;
		END IF;
	END IF;
END IF;
END PROCESS CONTADOR_DECADA;
END PROGRAMA;