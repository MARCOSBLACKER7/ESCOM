module boletaescom ( 
	clk,
	clr,
	en,
	display
	) ;

input  clk;
input  clr;
input  en;
inout [8:0] display;
