LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FFS IS 
	PORT(
		J, K, T, S, R, D: IN STD_LOGIC;
		CLK, CLR: IN STD_LOGIC;
		SEL: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		DISPLAY: OUT STD_LOGIC_VECTOR(5 DOWNTO O)
	);
ATTRIBUTE PIN_NUMBERS OF FFS: ENTITY IS
 " CLK:1 J:2 K:3 T:4 S:5 R:6 D:7 SEL(0):8 SEL(1):9" &
 " QJK:15 QSR:23 QT:14 QD:22 CLR:13 DISPLAY(0):16 DISPLAY(1):17 " &
 "DISPLAY(2):18 DISPLAY(3):19 DISPLAY(4):20 DISPLAY(5):21 " 
;
END FFS;

ARCHITECTURE PRACTICA OF FFS IS 
SIGNAL QJK:STD_LOGIC;
SIGNAL QSR:STD_LOGIC;
SIGNAL QT:STD_LOGIC;
SIGNAL QD:STD_LOGIC;

BEGIN 
	FFJK: PROCESS(CLK, CLR)
	BEGIN
	IF( CLR = '1') THEN 
			QJK <= '0';
	ELSIF( CLK'EVENT AND CLK='1') THEN
		QJK <= (J AND NOT QJK) + (NOT K AND QJK);
	END IF;
	END PROCESS FFJK;

	FFSR: PROCESS(CLK, CLR)
	BEGIN
	IF( CLR = '1') THEN 
			QSR <= '0';
	ELSIF( CLK'EVENT AND CLK='1') THEN
		QSR <= S + (NOT R AND  QRS);
	END IF;
	END PROCESS FFSR;

	FFT: PROCESS(CLK, CLR)
	BEGIN
	IF( CLR = '1') THEN 
			QT <= '0';
	ELSIF( CLK'EVENT AND CLK='1') THEN
		QT <= T XOR QT;
	END IF;
	END PROCESS FFT;

	FFD: PROCESS(CLK, CLR)
	BEGIN
	IF( CLR = '1') THEN 
			QD <= '0';
	ELSIF( CLK'EVENT AND CLK='1') THEN
		QT <= D;
	END IF;
	END PROCESS FFD;
	


	SELE: PROCESS(QJK, QSR, QT, QD, SEL)
	BEGIN 
   	IF QJK= '0' THEN DISPLAY <= "000000";
			ELSIF QJK= '1' THEN DISPLAY <= "100111";
			ELSIF QT= '0' THEN DISPLAY <= "000000";
			ELSIF QT= '1' THEN DISPLAY <= "100111";
			ELSIF QD= '0' THEN DISPLAY <= "000000";
			ELSIF QD= '1' THEN DISPLAY <= "100111";
			ELSIF QSR= '0' THEN DISPLAY <= "000000";
			ELSIF QSR= '1' THEN DISPLAY <= "100111";
		END IF 
		CASE SEL IS
		 WHEN "00" => DISPLAY <= QJK;
		 WHEN "01" => DISPLAY <= QT;
		 WHEN "10" => DISPLAY <= QD;
	     WHEN "11" => DISPLAY <= QSR;
		 WHEN OTHERS DISPLAY <= "ZZZZZZ";
		 END CASE;
	 END PROCESS SELE;



END PRACTICA;





