LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CONVERTIDOR IS
	PORT(
		CLK, CLR : IN STD_LOGIC;
		E0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		E1: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		DISPLAY: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		AN: INOUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);

	ATTRIBUTE PIN_NUMBERS OF CONVERTIDOR : ENTITY IS
		"CLK:1   "	    	&
		"CLR:13  "	    	&
		"E1(2):5 "		&
		"E1(1):6 "		&
		"E1(0):7 "		&
		"E0(3):8 "		&
		"E0(2):9 "		&
		"E0(1):10 "		&
		"E0(0):11 "     	&
		"AN(0):14 "     	&
		"AN(1):23 "     	&
		"AN(2):22 "     	&
		"DISPLAY(0):15 "   	&   
        "DISPLAY(1):16 "   	&   
       	"DISPLAY(2):17 "   	&  
 	    "DISPLAY(3):18 "   	&  
		"DISPLAY(4):19 "   	&  
		"DISPLAY(5):20 "   	&  
		"DISPLAY(6):21 ";   
END CONVERTIDOR;

ARCHITECTURE PROGRAMA OF CONVERTIDOR IS
CONSTANT CERO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0000001";
CONSTANT UNO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "1001111";
CONSTANT DOS : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0010010";
CONSTANT TRES : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0000110";
CONSTANT CUATRO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "1001100";
CONSTANT CINCO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0100100";
CONSTANT SEIS : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0100000";
CONSTANT SIETE : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0001111";
CONSTANT OCHO : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0000000";
CONSTANT NUEVE : STD_LOGIC_VECTOR(6 DOWNTO 0):=    "0000100";
CONSTANT BCDCERO : STD_LOGIC_VECTOR(3 DOWNTO 0):=   	 "0000";
CONSTANT BCDUNO : STD_LOGIC_VECTOR(3 DOWNTO 0):=    	 "0001";
CONSTANT BCDDOS : STD_LOGIC_VECTOR(3 DOWNTO 0):=   	 "0010";
CONSTANT BCDTRES : STD_LOGIC_VECTOR(3 DOWNTO 0):=   	 "0011";
CONSTANT BCDCUATRO : STD_LOGIC_VECTOR(3 DOWNTO 0):=    	 "0100";
CONSTANT BCDCINCO : STD_LOGIC_VECTOR(3 DOWNTO 0):=    	 "0101";
CONSTANT BCDSEIS : STD_LOGIC_VECTOR(3 DOWNTO 0):=    	 "0110";
CONSTANT BCDSIETE : STD_LOGIC_VECTOR(3 DOWNTO 0):=    	 "1011";
CONSTANT BCDOCHO : STD_LOGIC_VECTOR(3 DOWNTO 0):=    	 "1000";
CONSTANT BCDNUEVE : STD_LOGIC_VECTOR(3 DOWNTO 0):=    	 "1001";
SIGNAL BCD: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL E2:  STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	E2<=(OTHERS=>'0');
	ANILLO: PROCESS(CLK, CLR)
	BEGIN
		IF CLR = '1' THEN
			AN<="110";
		ELSIF RISING_EDGE(CLK) THEN
			AN<=TO_STDLOGICVECTOR(TO_BITVECTOR(AN) ROL 1);
		END IF;
	END PROCESS ANILLO;

	MUX: PROCESS(AN)
	BEGIN
		CASE AN IS
		WHEN "110"=>
			BCD<= E0;
		WHEN "101"=>
			BCD(3)<= '0';
			BCD(2)<= E1(2);
			BCD(1)<= E1(1);
			BCD(0)<= E1(0);
		WHEN "011"=>
			BCD<= E2;
		WHEN OTHERS =>
			BCD<=(OTHERS =>'-');
		END CASE;
	END PROCESS MUX;

	CO: PROCESS(BCD)
	BEGIN
		CASE BCD IS
		WHEN BCDCERO=>
			DISPLAY<= CERO;
		WHEN BCDUNO=>
			DISPLAY<= UNO;
		WHEN BCDDOS=>
			DISPLAY<= DOS;
		WHEN BCDTRES=>
			DISPLAY<= TRES;
		WHEN BCDCUATRO=>
			DISPLAY<= CUATRO;
		WHEN BCDCINCO=>
			DISPLAY<= CINCO;
		WHEN BCDSEIS=>
			DISPLAY<= SEIS;
		WHEN BCDSIETE=>
			DISPLAY<= SIETE;
		WHEN BCDOCHO=>
			DISPLAY<= OCHO;
		WHEN BCDNUEVE=>
			DISPLAY<= NUEVE;
		WHEN OTHERS =>
			DISPLAY<= (OTHERS =>'-');
		END CASE;
	END PROCESS CO;
END PROGRAMA;