module mensaje ( 
	clk,
	clr,
	an,
	d
	) ;

input  clk;
input  clr;
inout [2:0] an;
inout [6:0] d;
