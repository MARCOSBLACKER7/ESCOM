module secuencia ( 
	clk,
	clr,
	x,
	an0,
	d
	) ;

input  clk;
input  clr;
input  x;
inout  an0;
inout [6:0] d;
