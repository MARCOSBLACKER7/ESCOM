LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTADOR IS
	GENERIC( N : INTEGER := 4 );
	PORT(
		EN,CLR,CLK: IN STD_LOGIC;
		DISPLAY : INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);

	ATTRIBUTE PIN_NUMBERS OF CONTADOR: ENTITY IS 
        "CLK:1 "         &
        "CLR:13 "        &
        "EN:2 "          &
        "DISPLAY(0):15 " &
        "DISPLAY(1):16 " &
        "DISPLAY(2):17 " &
        "DISPLAY(3):18 " &
        "DISPLAY(4):19 " &
        "DISPLAY(5):20 " &
        "DISPLAY(6):21";
END CONTADOR;

ARCHITECTURE PROGRAMA OF CONTADOR IS
CONSTANT D0 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001111";
CONSTANT D1 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0010010";
CONSTANT D2 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000110";
CONSTANT D3 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001100";
CONSTANT D4 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100100";
CONSTANT D5 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100000";

BEGIN
	PCONT : PROCESS( CLK, CLR )
	BEGIN
		IF( CLR = '1' )THEN
			DISPLAY <= D0;
		ELSIF RISING_EDGE(CLK) THEN
		IF EN ='1' THEN
				IF DISPLAY = D0 THEN
					DISPLAY <= D1;
				ELSIF DISPLAY = D1 THEN
					DISPLAY <= D2;
				ELSIF DISPLAY = D2 THEN
					DISPLAY <= D3;
				ELSIF DISPLAY = D3 THEN
					DISPLAY <= D4;
				ELSIF DISPLAY = D4 THEN
					DISPLAY <= D5;

				ELSE
				DISPLAY<= D0;
				END IF;	
			END IF;
			END IF;
	END PROCESS PCONT;
END PROGRAMA;
