module numeros2 ( 
	en,
	clk,
	clr,
	upd,
	l,
	d,
	q,
	c
	) ;

input  en;
input  clk;
input  clr;
input  upd;
input  l;
input [6:0] d;
inout [6:0] q;
inout  c;
