library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CODIGO is
    Port ( BCD : in  STD_LOGIC_VECTOR (3 downto 0);
           DISPLAY : out  STD_LOGIC_VECTOR (6 downto 0));
end CODIGO;

architecture CONVERTIDOR of CODIGO is

begin


end CONVERTIDOR;

