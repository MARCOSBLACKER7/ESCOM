library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CONVERTIDOR is
    Port ( BCD : in  STD_LOGIC_VECTOR (3 downto 0);
           SEG : out  STD_LOGIC_VECTOR (6 downto 0));
end CONVERTIDOR;

architecture PROGRAMA of CONVERTIDOR is

--ABCDEFG	DIG
--0000001	0
--1001111	1
--0010010	2
--0000110	3
--1001100	4
--0100100	5
--0100000	6
--0001111	7
--0000000	8
--0000100	9

CONSTANT DIG0 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
CONSTANT DIG1 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
CONSTANT DIG2 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
CONSTANT DIG3 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
CONSTANT DIG4 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001100";
CONSTANT DIG5 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
CONSTANT DIG6 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100000";
CONSTANT DIG7 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001111";
CONSTANT DIG8 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
CONSTANT DIG9 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";

begin

	SEG <=	DIG0 WHEN ( BCD = X"0" ) ELSE
				DIG1 WHEN ( BCD = X"1" ) ELSE
				DIG2 WHEN ( BCD = X"2" ) ELSE
				DIG3 WHEN ( BCD = X"3" ) ELSE
				DIG4 WHEN ( BCD = X"4" ) ELSE
				DIG5 WHEN ( BCD = X"5" ) ELSE
				DIG6 WHEN ( BCD = X"6" ) ELSE
				DIG7 WHEN ( BCD = X"7" ) ELSE
				DIG8 WHEN ( BCD = X"8" ) ELSE
				DIG9; 
				
end PROGRAMA;
