LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REGISTRO IS 
	PORT(
		CLK, CLR, ES: IN STD_LOGIC;
		OPER: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	    D	: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		Q	: INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)

	);
ATTRIBUTE PIN_NUMBERS OF FFS: ENTITY IS
 
END REGISTRO;

ARCHITECTURE PRACTICA OF REGISTRO IS 
BEGIN
	PREG : PROCESS (CLR, CLK)
	BEGIN
		IF(CLR= '1') THEN
			Q<= (OTHERS =>  '0');	--Q<= "0000"; --Q <= X"0";
		ELSIF(CLK EVENT AND CLK = '1' ) THEN
		
		FOR I IN  3 DOWNTO 0 LOOP
			IF(I = 0 ) THEN

		 	Q(I)<=  ( Q(I)   AND NOT OPER(1) AND NOT OPER(0) ) OR
					( D(I)   AND NOT OPER(1) AND     OPER(0) ) OR
					( ES     AND     OPER(1) AND NOT OPER(0) ) OR
					( Q(I+1) AND     OPER(1) AND     OPER(0) );
			
			ELSIF (I = 3) THEN
			Q(I)<=  ( Q(I)   AND NOT OPER(1) AND NOT OPER(0) ) OR
					( D(I)   AND NOT OPER(1) AND     OPER(0) ) OR
					(Q(I-1)  AND     OPER(1) AND NOT OPER(0) ) OR
					(ES      AND     OPER(1) AND     OPER(0) );


			ELSE

	Q(I)<=  ( Q(I) AND NOT OPER(1) AND NOT OPER(0) ) OR
			( D(I) AND NOT OPER(1) AND     OPER(0) ) OR
			( Q(I-1) AND     OPER(1) AND NOT OPER(0) ) OR
			( Q(I+1)   AND     OPER(1) AND     OPER(0) );
			END LOOP;
			END IF;
 	END PROCESS PREG;
END PRACTICA;





