LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FFL IS
	PORT( J, K, T, D, S, R: IN STD_LOGIC;
		  CLK, CLR: IN STD_LOGIC;
		  SEL: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		  DISPLAY: OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
		);

	ATTRIBUTE PIN_NUMBERS OF FFL: ENTITY IS
		"DISPLAY(0):16 DISPLAY(1):17 DISPLAY(2):18"
		& " DISPLAY(3):19 DISPLAY(4):20 DISPLAY(5):21"
		& " CLK:1 CLR:13 J:2 K:3 T:4 S:5 R:6 D:7"
		& " SEL(0):8 SEL(1):9";
END FFL;

ARCHITECTURE FFS OF FFL IS
	SIGNAL QJK, QD, QT, QSR, Q: STD_LOGIC;
	
	BEGIN
		FFJK: PROCESS(CLK,CLR)
		BEGIN
			IF (CLR='1') THEN
				QJK <= '0';
			ELSIF(CLK'EVENT AND CLK='1') THEN
				QJK <= (J AND (NOT QJK))OR((NOT K) AND QJK);
			END IF;
		END PROCESS FFJK;

		FFD: PROCESS(CLK,CLR)
		BEGIN
			IF (CLR='1') THEN
				QD <= '0';
			ELSIF(CLK'EVENT AND CLK='1') THEN
				QD <= D;
			END IF;
		END PROCESS FFD;
		

		FFT: PROCESS(CLK,CLR)
		BEGIN
			IF (CLR='1') THEN
				QT <= '0';
			ELSIF(CLK'EVENT AND CLK='1') THEN
				QT <= T XOR QT;
			END IF;
		END PROCESS FFT;

		FFSR: PROCESS(CLK,CLR)
		BEGIN
			IF (CLR='1') THEN
				QSR <= '0';
			ELSIF(CLK'EVENT AND CLK='1') THEN
				QSR <= S OR ((NOT R) AND QSR);
			END IF;
		END PROCESS FFSR;

		WITH SEL SELECT 
		Q <= QJK WHEN "00",
			 QT WHEN "01",
			 QD WHEN "10",
			 QSR WHEN OTHERS;

		DISPLAY <= 	"000000" WHEN( Q = '0' )ELSE 
					"100111";
END FFS;
