LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REGISTRO IS 
	PORT(
		CLK, CLR, ES: IN STD_LOGIC;
		OPER: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	    D	: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		Q	: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0)

	);
ATTRIBUTE PIN_NUMBERS OF FFS: ENTITY IS
 
END REGISTRO;

ARCHITECTURE PRACTICA OF REGISTRO IS 
BEGIN
	PREG : PROCESS (CLR, CLK)
	BEGIN
		IF(CLR= '1') THEN
			Q<= (OTHERS =>  '0');	--Q<= "0000"; --Q <= X"0";
		ELSIF(CLK EVENT AND CLK = '1' ) THEN

 	Q(0)<=  ( Q(0) AND NOT OPER(1) AND NOT OPER(0) ) OR
			( D(0) AND NOT OPER(1) AND     OPER(0) ) OR
			( ES   AND     OPER(1) AND NOT OPER(0) ) OR
			( Q(1) AND     OPER(1) AND     OPER(0) );

	Q(1)<=  ( Q(1) AND NOT OPER(1) AND NOT OPER(0) ) OR
			( D(1) AND NOT OPER(1) AND     OPER(0) ) OR
			( Q(0) AND     OPER(1) AND NOT OPER(0) ) OR
			( Q(2) AND     OPER(1) AND     OPER(0) );

	Q(2)<=  ( Q(2) AND NOT OPER(1) AND NOT OPER(0) ) OR
			( D(2) AND NOT OPER(1) AND     OPER(0) ) OR
			( Q(1) AND     OPER(1) AND NOT OPER(0) ) OR
			( Q(3) AND     OPER(1) AND     OPER(0) );

	Q(3)<=  ( Q(3) AND NOT OPER(1) AND NOT OPER(0) ) OR
			( D(3) AND NOT OPER(1) AND     OPER(0) ) OR
			( Q(2) AND     OPER(1) AND NOT OPER(0) ) OR
			( ES   AND     OPER(1) AND     OPER(0) );
		END IF;
 	END PROCESS PREG;
END PRACTICA;





