module numeros ( 
	en,
	clk,
	clr,
	q
	) ;

input  en;
input  clk;
input  clr;
inout [6:0] q;
