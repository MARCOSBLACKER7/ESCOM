module sincrono ( 
	clk,
	clr,
	e,
	d1,
	d2,
	uni,
	dec
	) ;

input  clk;
input  clr;
inout  e;
inout  d1;
inout  d2;
inout [3:0] uni;
inout [2:0] dec;
