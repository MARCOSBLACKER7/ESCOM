LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY HEXADECIMAL IS
	PORT(
		CLK, CLR, EN : IN STD_LOGIC;
		DISPLAY : INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
ATTRIBUTE PIN_NUMBERS OF HEXADECIMAL: ENTITY IS 
        "CLK:1 "         &
        "CLR:13 "        &
        "EN:2 "          &
        "DISPLAY(0):15 " &
        "DISPLAY(1):16 " &
        "DISPLAY(2):17 " &
        "DISPLAY(3):18 " &
        "DISPLAY(4):19 " &
        "DISPLAY(5):20 " &
        "DISPLAY(6):21";

END HEXADECIMAL;

ARCHITECTURE PROGRAMA OF HEXADECIMAL IS
CONSTANT Q0  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
CONSTANT Q1  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
CONSTANT Q2  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
CONSTANT Q3  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
CONSTANT Q4  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001100";
CONSTANT Q5  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
CONSTANT Q6  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100000";
CONSTANT Q7  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001111";
CONSTANT Q8  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
CONSTANT Q9  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";
CONSTANT Q10 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001000";
CONSTANT Q11 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1100000";
CONSTANT Q12 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110001";
CONSTANT Q13 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1000010";
CONSTANT Q14 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000";
CONSTANT Q15 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0111000";

BEGIN
PMSJ : PROCESS(CLK, CLR)
BEGIN
IF(CLR = '1') THEN
  DISPLAY <= Q0;
	ELSIF RISING_EDGE(CLK) THEN
        IF EN = '1' THEN
            IF DISPLAY = Q0 THEN
                DISPLAY <= Q1;
            ELSIF DISPLAY = Q1 THEN
                DISPLAY <= Q2;
            ELSIF DISPLAY = Q2 THEN
                DISPLAY <= Q3;
            ELSIF DISPLAY = Q3 THEN
                DISPLAY <= Q4;
            ELSIF DISPLAY = Q4 THEN
                DISPLAY <= Q5;
            ELSIF DISPLAY = Q5 THEN
                DISPLAY <= Q6;
            ELSIF DISPLAY = Q6 THEN
                DISPLAY <= Q7;
            ELSIF DISPLAY = Q7 THEN
                DISPLAY <= Q8;
            ELSIF DISPLAY = Q8 THEN
                DISPLAY <= Q9;
            ELSIF DISPLAY = Q9 THEN
                DISPLAY <= Q10;
            ELSIF DISPLAY = Q10 THEN
                DISPLAY <= Q11;
            ELSIF DISPLAY = Q11 THEN
                DISPLAY <= Q12;
            ELSIF DISPLAY = Q12 THEN
                DISPLAY <= Q13;
            ELSIF DISPLAY = Q13 THEN
                DISPLAY <= Q14;
            ELSIF DISPLAY = Q14 THEN
                DISPLAY <= Q15;
                
            ELSE
                DISPLAY <= Q0;
            END IF;
        END IF;
	END IF;
END PROCESS PMSJ;
END PROGRAMA;
