LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY BOLETAESCOM IS
	PORT(
		CLK, CLR, EN : IN STD_LOGIC;
		DISPLAY : INOUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
ATTRIBUTE PIN_NUMBERS OF BOLETAESCOM : ENTITY IS
        "CLK:1 "         &
        "CLR:13 "        &
        "EN:2 "          &
        "DISPLAY(0):15 " &
        "DISPLAY(1):16 " &
        "DISPLAY(2):17 " &
        "DISPLAY(3):18 " &
        "DISPLAY(4):19 " &
        "DISPLAY(5):20 " &
        "DISPLAY(6):21";

END BOLETAESCOM;

ARCHITECTURE PROGRAMA OF BOLETAESCOM IS
--2016601777
CONSTANT CERO :   STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
CONSTANT UNO:     STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
CONSTANT DOS :    STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
CONSTANT TRES :   STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
CONSTANT CUATRO : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001100";
CONSTANT CINCO :  STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
CONSTANT SEIS :   STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100000";
CONSTANT SIETE :  STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001111";
CONSTANT OCHO :   STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
CONSTANT NUEVE :  STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";

CONSTANT ETI00 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
CONSTANT ETI01 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
CONSTANT ETI10 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";

CONSTANT Q0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & DOS;  
CONSTANT Q1 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & CERO;
CONSTANT Q2 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & UNO;
CONSTANT Q3 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & SEIS;
CONSTANT Q4 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI01 & SEIS;
CONSTANT Q5 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI01 & CERO;
CONSTANT Q6 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI01 & UNO;
CONSTANT Q7 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & SIETE;
CONSTANT Q8 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI01 & SIETE;
CONSTANT Q9 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI10 & SIETE;

BEGIN
PMSJ : PROCESS(CLK, CLR)
BEGIN
IF(CLR = '1') THEN
	DISPLAY <= Q0;
	ELSIF RISING_EDGE(CLK) THEN
        IF EN = '1' THEN
            IF DISPLAY = Q0 THEN
                DISPLAY <= Q1;
            ELSIF DISPLAY = Q1 THEN
                DISPLAY <= Q2;
            ELSIF DISPLAY = Q2 THEN
                DISPLAY <= Q3;
            ELSIF DISPLAY = Q3 THEN
                DISPLAY <= Q4;
            ELSIF DISPLAY = Q4 THEN
                DISPLAY <= Q5;
            ELSIF DISPLAY = Q5 THEN
                DISPLAY <= Q6;
            ELSIF DISPLAY = Q6 THEN
                DISPLAY <= Q7;
            ELSIF DISPLAY = Q7 THEN
                DISPLAY <= Q8;
            ELSIF DISPLAY = Q8 THEN
                DISPLAY <= Q9;
                
            ELSE
                DISPLAY <= Q0;
                END IF;
            END IF;
	END IF;
END PROCESS PMSJ;
END PROGRAMA;
