library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BCD27SEG is
    Port ( BCD : in  STD_LOGIC_VECTOR (3 downto 0);
           SEG : out  STD_LOGIC_VECTOR (6 downto 0));
end BCD27SEG;

architecture PROGRAMA of BCD27SEG is
CONSTANT DIG0 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
CONSTANT DIG1 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
CONSTANT DIG2 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
CONSTANT DIG3 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
CONSTANT DIG4 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001100";
CONSTANT DIG5 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
CONSTANT DIG6 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100000";
CONSTANT DIG7 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001110";
CONSTANT DIG8 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
CONSTANT DIG9 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";

begin
		SEG <= DIG0 WHEN (BCD = "0000" ) ELSE
				 DIG1 WHEN (BCD = "0001" ) ELSE
				 DIG2 WHEN (BCD = "0010" ) ELSE
				 DIG3 WHEN (BCD = "0011" ) ELSE
				 DIG4 WHEN (BCD = "0100" ) ELSE
				 DIG5 WHEN (BCD = "0101" ) ELSE
				 DIG6 WHEN (BCD = "0110" ) ELSE
				 DIG7 WHEN (BCD = "0111" ) ELSE
				 DIG8 WHEN (BCD = "1000" ) ELSE
				 DIG9 WHEN (BCD = "1001" ) ELSE
 				 "1111111";
				 

end PROGRAMA;

