LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MSJ IS
	PORT(
		CLK, CLR, EN : IN STD_LOGIC;
		DISPLAY : INOUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
ATTRIBUTE PIN_NUMBERS OF MSJ: ENTITY IS 
        "CLK:1 "         &
        "CLR:13 "        &
        "EN:2 "          &
        "DISPLAY(0):15 " &
        "DISPLAY(1):16 " &
        "DISPLAY(2):17 " &
        "DISPLAY(3):18 " &
        "DISPLAY(4):19 " &
        "DISPLAY(5):20 " &
        "DISPLAY(6):21";

END MSJ;

ARCHITECTURE PROGRAMA OF MSJ IS
CONSTANT Ld : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1000010";
CONSTANT LI : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
CONSTANT LS : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
CONSTANT LE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000";
CONSTANT Ln : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0101010";
CONSTANT LO : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
CONSTANT LG : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";
CONSTANT LT : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110000";
CONSTANT LA : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001000";
CONSTANT LL : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110001";

CONSTANT ETI00 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
CONSTANT ETI01 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
CONSTANT ETI10 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";

CONSTANT Q0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & Ld;
CONSTANT Q1 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & LI;
CONSTANT Q2 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & LS;
CONSTANT Q3 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & LE;
CONSTANT Q4 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & Ln;
CONSTANT Q5 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & LO;
CONSTANT Q6 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI01 & Ld;
CONSTANT Q7 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI01 & LI;
CONSTANT Q8 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & LG;
CONSTANT Q9 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI10 & LI;
CONSTANT Q10 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & LT;
CONSTANT Q11 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & LA;
CONSTANT Q12 : STD_LOGIC_VECTOR(8 DOWNTO 0) := ETI00 & LL;

BEGIN
	PMSJ : PROCESS(CLK, CLR)
	BEGIN
		IF(CLR = '1') THEN
		  DISPLAY <= q0;
		  ELSIF RISING_EDGE(CLK) THEN
                IF EN = '1' THEN
                    IF DISPLAY = Q0 THEN
                        DISPLAY <= Q1;
                    ELSIF DISPLAY = Q1 THEN
                        DISPLAY <= Q2;
                    ELSIF DISPLAY = Q2 THEN
                        DISPLAY <= Q3;
                    ELSIF DISPLAY = Q3 THEN
                        DISPLAY <= Q4;
                    ELSIF DISPLAY = Q4 THEN
                        DISPLAY <= Q5;
                    ELSIF DISPLAY = Q5 THEN
                        DISPLAY <= Q6;
                    ELSIF DISPLAY = Q6 THEN
                        DISPLAY <= Q7;
                    ELSIF DISPLAY = Q7 THEN
                        DISPLAY <= Q8;
                    ELSIF DISPLAY = Q8 THEN
                        DISPLAY <= Q9;
                    ELSIF DISPLAY = Q9 THEN
                        DISPLAY <= Q10;
                    ELSIF DISPLAY = Q10 THEN
                        DISPLAY <= Q11;
                    ELSIF DISPLAY = Q11 THEN
                        DISPLAY <= Q12;

                    ELSE
                        DISPLAY <= Q0;
                    END IF;
	           END IF;
			END IF;
	END PROCESS PMSJ;
END PROGRAMA;
